/**
 * Testbench:
 *  bias_add
 *
 * Created:
 *  Fri Jan 10 21:56:05 AEDT 2020
 *
 * Author:
 *  Berin Martini (berin.martini@gmail.com)
 */

`timescale 1ns/10ps

`define TB_VERBOSE
//`define VERBOSE


`include "bias_add.sv"

module bias_add_tb;

    /**
     * Clock and control functions
     */

    // Generate a clk
    reg clk = 0;
    always #1 clk = !clk;

    // End of simulation event definition
    event end_trigger;
    always @(end_trigger) $finish;

`ifdef TB_VERBOSE
    // Display header information
    initial #1 display_header();
    always @(end_trigger) display_header();

    // And strobe signals at each clk
    always @(posedge clk) display_signals();
`endif

//    initial begin
//        $dumpfile("result.vcd"); // Waveform file
//        $dumpvars;
//    end


    /**
     * Local parameters
     */

    localparam NUM_WIDTH    = 16;
    localparam NUM_POINT    = 8;


    // transform signed fixed point representation to real
    function real num_f2r;
        input signed [NUM_WIDTH-1:0] value;

        begin
            num_f2r = value / ((1<<NUM_POINT) * 1.0);
        end
    endfunction

    // transform real to signed fixed point representation
    function signed [NUM_WIDTH-1:0] num_r2f;
        input real value;

        begin
            num_r2f = value * (1<<(NUM_POINT));
        end
    endfunction


`ifdef TB_VERBOSE
    initial begin
        $display("Testbench for 'bias_add'");
    end
`endif


    /**
     *  signals, registers and wires
     */

    reg         [NUM_WIDTH-1:0] bias;
    reg         [NUM_WIDTH-1:0] up_data;
    wire signed [NUM_WIDTH-1:0] dn_data;


    reg                         up_valid;
    reg                         dn_valid;


    /**
     * Unit under test
     */

    bias_add #(
        .NUM_WIDTH  (NUM_WIDTH))
    uut (
        .clk        (clk),

        .bias       (bias),

        .up_data    (up_data),
        .dn_data    (dn_data)
    );


    // one pipeline depth
    always @(posedge clk)
        dn_valid <= up_valid;


    /**
     * Wave form display
     */

    task display_signals;
        $display(
            "%d",
            $time,

            "\t<bias> %f",
            num_f2r(bias),

            "\t<up> %b %f  ",
            up_valid,
            num_f2r(up_data),

            "\t<dn> %b %f",
            dn_valid,
            num_f2r(dn_data),

        );

    endtask // display_signals

    task display_header;
        $display(
            "\t\ttime",

            "\t\tbias",

            "\t\tup",

            "\t\t\tdn",
        );
    endtask


    /**
     * Testbench program
     */

    initial begin
        // init values

        bias        = num_r2f(2.5);
        up_data     = 'b0;
        up_valid    = 1'b0;

        //end init

        repeat(5) @(negedge clk);

`ifdef TB_VERBOSE
    $display("send data");
`endif
        @(negedge clk);

        repeat(20) begin
            up_valid    <= 1'b1;
            up_data     <= num_r2f(num_f2r(up_data)+1.0);
            @(negedge clk);
        end

        up_valid    <= 1'b0;
        up_data     <= 'b0;
        repeat(10) @(negedge clk);


`ifdef TB_VERBOSE
    $display("END");
`endif
        -> end_trigger;
    end

endmodule
