    localparam
        CFG_LAYERS   =  0,
        CFG_KER_WR   =  1,
        CFG_KER_RD   =  2;
