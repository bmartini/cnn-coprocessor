    localparam
        CFG_LAYERS       =  0,
        CFG_KER_WR       =  1,
        CFG_KER_RD       =  2,
        CFG_IMG_WR       =  3,
        CFG_IMG_RD       =  4,
        CFG_IR_IMG_W     =  5,
        CFG_IR_IMG_DH    =  6,
        CFG_IR_PAD       =  7,
        CFG_IR_CONV      =  8,
        CFG_IW_IMG_W     =  9,
        CFG_IW_START     = 10,
        CFG_IW_STEP      = 11;
