    localparam
        CFG_LAYERS   =  0;
